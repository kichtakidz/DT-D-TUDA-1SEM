`timescale 1ns / 1ns

module s_box_1

    ( input   logic [3:0] I,  // 4-bit input
      output  logic [3:0] O); // substituted output

/* ====================================== INSERT CODE HERE ====================================== */
  


/* ============================================================================================== */

endmodule