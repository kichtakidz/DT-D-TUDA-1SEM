`timescale 1ns / 1ns

module p_box

    ( input   logic [7:0] I,   // 8-bit input
      output  logic [7:0] O); // rearranged output

/* ====================================== INSERT CODE HERE ====================================== */



/* ============================================================================================== */

endmodule

