`timescale 1ns / 1ns

module key_schedule

    ( input   logic [31:0] K,               // 32-bit key
      output  logic [7:0] K0, K1, K2, K3);  // round keys

/* ====================================== INSERT CODE HERE ====================================== */
 

 
/* ============================================================================================== */

endmodule
